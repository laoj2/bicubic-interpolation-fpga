library verilog;
use verilog.vl_types.all;
entity tb_c_unit is
end tb_c_unit;
